`ifndef __CRYPTO_DPI_TESTS_SV__
`define __CRYPTO_DPI_TESTS_SV__

`include "tests/crypto_dpi_aes_ecb_test.sv"
`include "tests/crypto_dpi_evp_test.sv"

`endif
